module top(
input [3:0] A,
input [3:0] B,
input [2:0] ALUctr,
output reg [3:0] ALUout,
output reg [3:0] temp,
output reg less,
output reg of,zf,cf

);

always@(*)begin
	ALUout = 4'b0;



end


endmodule
