module top(
	input clk,
	input rst,
	output a
);




endmodule
